////////////////////////////////////////////////////////////////////////////////
// @file    tb_top_axis.v
// @author  JAY CONVERTINO
// @date    2022.10.24
// @brief   Generic AXIS test bench top with verification.
// @details This generic top and mod axis test bench is created for a FIFO.
//          It will have to be altered for other devices that alter the input
//          for some sort of output.
////////////////////////////////////////////////////////////////////////////////

`timescale 1 ns/10 ps

module tb_axis;
  //parameter or local param bus, user and dest width? and files as well? 
  
  localparam CLK_PERIOD = 500;
  localparam RST_PERIOD = 1000;
  
  wire        tb_m_clk;
  wire        tb_m_rstn;
  wire        tb_dut_valid;
  wire        tb_dut_ready;
  wire        tb_dut_data;
  wire        tb_dut_keep;
  wire        tb_dut_last;
  wire        tb_dut_user;
  wire        tb_dut_dest;
  
  wire        tb_s_clk;
  wire        tb_s_rstn;
  wire        tb_stim_valid;
  wire        tb_stim_data;
  wire        tb_stim_keep;
  wire        tb_stim_last;
  wire        tb_stim_user;
  wire        tb_stim_dest;
  
  reg         tb_cnt_clk  = 0;
  reg         tb_cnt_rstn = 0;
  wire        tb_cnt_data;
  
  clk_stimulator #(
    .CLOCKS(2), // # of clocks
    .CLOCK_BASE(1000000), // clock time base mhz
    .CLOCK_DIFFS(100), // clock time diff mhz
    .RESETS(2), // # of resets
    .RESET_BASE(200), // time to stay in reset
    .RESET_DIFFS(100) // time diff for other resets
  ) clk_stim
  (
    //clk out ... maybe a vector of clks with diff speeds.
    .clkv(tb_dut_clk, tb_stim_clk),
    //rstn out ... maybe a vector of rsts with different off times
    .rstnv(tb_dut_rstn, tb_stim_rstn),
    .rstv()
  );
  
  
  axis_stimulator #(
    .BUS_WIDTH(1),
    .USER_WIDTH(1),
    .DEST_WIDTH(1),
    .FILE_IN(),
    .FILE_OUT()
  ) axis_stim
  (
    // read
    .m_axis_aclk(tb_stim_clk),
    .m_axis_arstn(tb_stim_rstn),
    .m_axis_tvalid(tb_stim_valid),
    .m_axis_tready(tb_stim_ready),
    .m_axis_tdata(tb_stim_data),
    .m_axis_tkeep(tb_stim_keep),
    .m_axis_tlast(tb_stim_last),
    .m_axis_tuser(tb_stim_user),
    .m_axis_tdest(tb_stim_dest),
    // write
    .s_axis_aclk(tb_dut_clk),
    .s_axis_arstn(tb_dut_rstn),
    .s_axis_tvalid(tb_dut_valid),
    .s_axis_tready(tb_dut_ready),
    .s_axis_tdata(tb_dut_data),
    .s_axis_tkeep(tb_dut_keep),
    .s_axis_tlast(tb_dut_last),
    .s_axis_tuser(tb_dut_user),
    .s_axis_tdest(tb_dut_dest)
  );
  
  axis_fifo #(
    .FIFO_DEPTH(256),
    .COUNT_WIDTH(8),
    .BUS_WIDTH(1),
    .USER_WIDTH(1),
    .DEST_WIDTH(1),
    .RAM_TYPE("block"),
    .PACKET_MODE(0),
    .COUNT_DELAY(1),
    .COUNT_ENA(1)
  ) dut
  (
    // read
    .m_axis_aclk(tb_m_clk),
    .m_axis_arstn(tb_m_rstn),
    .m_axis_tvalid(tb_dut_valid),
    .m_axis_tready(tb_dut_ready),
    .m_axis_tdata(tb_dut_data),
    .m_axis_tkeep(tb_dut_keep),
    .m_axis_tlast(tb_dut_last),
    .m_axis_tuser(tb_dut_user),
    .m_axis_tdest(tb_dut_dest),
    // write
    .s_axis_aclk(tb_stim_clk),
    .s_axis_arstn(tb_stim_rstn),
    .s_axis_tvalid(tb_stim_valid),
    .s_axis_tready(tb_stim_ready),
    .s_axis_tdata(tb_stim_data),
    .s_axis_tkeep(tb_stim_keep),
    .s_axis_tlast(tb_stim_last),
    .s_axis_tuser(tb_stim_user),
    .s_axis_tdest(tb_stim_dest),
    // data count
    .data_count_aclk(tb_cnt_clk),
    .data_count_arstn(tb_cnt_rstn),
    .data_count(tb_cnt_data)
  );
    
endmodule

